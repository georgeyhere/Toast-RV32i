`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/04/2021 08:21:50 PM
// Design Name: 
// Module Name: toast_OOP_package
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


package toast_OOP_package;

    typedef enum int unsigned {inst_NOP = 0,
                               inst_LUI = 1} instruction_t;
    
    

endpackage
