@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00 
13 00 00 00 13 00 00 00 13 00 00 00 6F 00 C0 04 
73 2F 20 34 93 0F 80 00 63 0A FF 03 93 0F 90 00 
63 06 FF 03 93 0F B0 00 63 02 FF 03 17 0F 00 00 
13 0F 0F 00 63 04 0F 00 67 00 0F 00 73 2F 20 34 
63 54 0F 00 6F 00 40 00 93 E1 91 53 17 0F 00 00 
23 20 3F 00 6F F0 9F FF 93 00 00 00 13 01 00 00 
93 01 00 00 13 02 00 00 93 02 00 00 13 03 00 00 
93 03 00 00 13 04 00 00 93 04 00 00 13 05 00 00 
93 05 00 00 13 06 00 00 93 06 00 00 13 07 00 00 
93 07 00 00 13 08 00 00 93 08 00 00 13 09 00 00 
93 09 00 00 13 0A 00 00 93 0A 00 00 13 0B 00 00 
93 0B 00 00 13 0C 00 00 93 0C 00 00 13 0D 00 00 
93 0D 00 00 13 0E 00 00 93 0E 00 00 13 0F 00 00 
93 0F 00 00 73 25 40 F1 63 10 05 00 97 02 00 00 
93 82 02 00 73 90 52 30 73 50 00 18 97 02 00 00 
93 82 02 00 73 90 52 30 B7 02 00 80 93 82 F2 FF 
73 90 02 3B 93 02 F0 01 73 90 02 3A 73 50 40 30 
97 02 00 00 93 82 02 00 73 90 52 30 73 50 20 30 
73 50 30 30 93 01 00 00 97 02 00 00 93 82 02 00 
73 90 52 30 13 05 10 00 13 15 F5 01 63 4C 05 00 
0F 00 F0 0F 93 01 10 00 93 08 D0 05 13 05 00 00 
73 00 00 00 97 02 00 00 93 82 02 00 63 8A 02 00 
73 90 52 10 B7 B2 00 00 93 82 92 10 73 90 22 30 
73 50 00 30 97 02 00 00 93 82 02 00 73 90 12 34 
73 25 40 F1 73 00 20 30 93 00 00 00 13 01 00 00 
33 87 20 00 93 03 00 00 93 01 20 00 63 16 77 4C 
93 00 10 00 13 01 10 00 33 87 20 00 93 03 20 00 
93 01 30 00 63 1A 77 4A 93 00 30 00 13 01 70 00 
33 87 20 00 93 03 A0 00 93 01 40 00 63 1E 77 48 
93 00 00 00 37 81 FF FF 33 87 20 00 B7 83 FF FF 
93 01 50 00 63 12 77 48 B7 00 00 80 13 01 00 00 
33 87 20 00 B7 03 00 80 93 01 60 00 63 16 77 46 
B7 00 00 80 37 81 FF FF 33 87 20 00 B7 83 FF 7F 
93 01 70 00 63 1A 77 44 93 00 00 00 37 81 00 00 
13 01 F1 FF 33 87 20 00 B7 83 00 00 93 83 F3 FF 
93 01 80 00 63 1A 77 42 B7 00 00 80 93 80 F0 FF 
13 01 00 00 33 87 20 00 B7 03 00 80 93 83 F3 FF 
93 01 90 00 63 1A 77 40 B7 00 00 80 93 80 F0 FF 
37 81 00 00 13 01 F1 FF 33 87 20 00 B7 83 00 80 
93 83 E3 FF 93 01 A0 00 63 18 77 3E B7 00 00 80 
37 81 00 00 13 01 F1 FF 33 87 20 00 B7 83 00 80 
93 83 F3 FF 93 01 B0 00 63 18 77 3C B7 00 00 80 
93 80 F0 FF 37 81 FF FF 33 87 20 00 B7 83 FF 7F 
93 83 F3 FF 93 01 C0 00 63 18 77 3A 93 00 00 00 
13 01 F0 FF 33 87 20 00 93 03 F0 FF 93 01 D0 00 
63 1C 77 38 93 00 F0 FF 13 01 10 00 33 87 20 00 
93 03 00 00 93 01 E0 00 63 10 77 38 93 00 F0 FF 
13 01 F0 FF 33 87 20 00 93 03 E0 FF 93 01 F0 00 
63 14 77 36 93 00 10 00 37 01 00 80 13 01 F1 FF 
33 87 20 00 B7 03 00 80 93 01 00 01 63 16 77 34 
93 00 D0 00 13 01 B0 00 B3 80 20 00 93 03 80 01 
93 01 10 01 63 9A 70 32 93 00 E0 00 13 01 B0 00 
33 81 20 00 93 03 90 01 93 01 20 01 63 1E 71 30 
93 00 D0 00 B3 80 10 00 93 03 A0 01 93 01 30 01 
63 94 70 30 13 02 00 00 93 00 D0 00 13 01 B0 00 
33 87 20 00 13 03 07 00 13 02 12 00 93 02 20 00 
E3 14 52 FE 93 03 80 01 93 01 40 01 63 1E 73 2C 
13 02 00 00 93 00 E0 00 13 01 B0 00 33 87 20 00 
13 00 00 00 13 03 07 00 13 02 12 00 93 02 20 00 
E3 12 52 FE 93 03 90 01 93 01 50 01 63 16 73 2A 
13 02 00 00 93 00 F0 00 13 01 B0 00 33 87 20 00 
13 00 00 00 13 00 00 00 13 03 07 00 13 02 12 00 
93 02 20 00 E3 10 52 FE 93 03 A0 01 93 01 60 01 
63 1C 73 26 13 02 00 00 93 00 D0 00 13 01 B0 00 
33 87 20 00 13 02 12 00 93 02 20 00 E3 16 52 FE 
93 03 80 01 93 01 70 01 63 18 77 24 13 02 00 00 
93 00 E0 00 13 01 B0 00 13 00 00 00 33 87 20 00 
13 02 12 00 93 02 20 00 E3 14 52 FE 93 03 90 01 
93 01 80 01 63 12 77 22 13 02 00 00 93 00 F0 00 
13 01 B0 00 13 00 00 00 13 00 00 00 33 87 20 00 
13 02 12 00 93 02 20 00 E3 12 52 FE 93 03 A0 01 
93 01 90 01 63 1A 77 1E 13 02 00 00 93 00 D0 00 
13 00 00 00 13 01 B0 00 33 87 20 00 13 02 12 00 
93 02 20 00 E3 14 52 FE 93 03 80 01 93 01 A0 01 
63 14 77 1C 13 02 00 00 93 00 E0 00 13 00 00 00 
13 01 B0 00 13 00 00 00 33 87 20 00 13 02 12 00 
93 02 20 00 E3 12 52 FE 93 03 90 01 93 01 B0 01 
63 1C 77 18 13 02 00 00 93 00 F0 00 13 00 00 00 
13 00 00 00 13 01 B0 00 33 87 20 00 13 02 12 00 
93 02 20 00 E3 12 52 FE 93 03 A0 01 93 01 C0 01 
63 14 77 16 13 02 00 00 13 01 B0 00 93 00 D0 00 
33 87 20 00 13 02 12 00 93 02 20 00 E3 16 52 FE 
93 03 80 01 93 01 D0 01 63 10 77 14 13 02 00 00 
13 01 B0 00 93 00 E0 00 13 00 00 00 33 87 20 00 
13 02 12 00 93 02 20 00 E3 14 52 FE 93 03 90 01 
93 01 E0 01 63 1A 77 10 13 02 00 00 13 01 B0 00 
93 00 F0 00 13 00 00 00 13 00 00 00 33 87 20 00 
13 02 12 00 93 02 20 00 E3 12 52 FE 93 03 A0 01 
93 01 F0 01 63 12 77 0E 13 02 00 00 13 01 B0 00 
13 00 00 00 93 00 D0 00 33 87 20 00 13 02 12 00 
93 02 20 00 E3 14 52 FE 93 03 80 01 93 01 00 02 
63 1C 77 0A 13 02 00 00 13 01 B0 00 13 00 00 00 
93 00 E0 00 13 00 00 00 33 87 20 00 13 02 12 00 
93 02 20 00 E3 12 52 FE 93 03 90 01 93 01 10 02 
63 14 77 08 13 02 00 00 13 01 B0 00 13 00 00 00 
13 00 00 00 93 00 F0 00 33 87 20 00 13 02 12 00 
93 02 20 00 E3 12 52 FE 93 03 A0 01 93 01 20 02 
63 1C 77 04 93 00 F0 00 33 01 10 00 93 03 F0 00 
93 01 30 02 63 12 71 04 93 00 00 02 33 81 00 00 
93 03 00 02 93 01 40 02 63 18 71 02 B3 00 00 00 
93 03 00 00 93 01 50 02 63 90 70 02 93 00 00 01 
13 01 E0 01 33 80 20 00 93 03 00 00 93 01 60 02 
63 14 70 00 63 10 30 02 0F 00 F0 0F 63 80 01 00 
93 91 11 00 93 E1 11 00 93 08 D0 05 13 85 01 00 
73 00 00 00 0F 00 F0 0F 93 01 10 00 93 08 D0 05 
13 05 00 00 73 00 00 00 73 10 00 C0 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
@00000000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 
